module uart_retrans_fsm (
    input clk,
    input reset,
    input ack,
    input frame_valid,
    input parity_error,
    input timeout,
    output error,
    output request_resend,
    output valid);

    
    
endmodule
