module elc_top(
        input clk,
        input reset,
        input [2:0] in,
        input card_is_in,
        input enter,
        output unlock,
        output error,
        output card_is_needed);

        

endmodule
