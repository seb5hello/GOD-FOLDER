module elc #(parameter [2:0] code = 3'b000)(
        input clk,
        input reset,
        input [2:0] in,
        input card_is_in,
        input enter,
        input tL,
        input tS,
        output trL,
        output trS,
        output unlock,
        output error,
        output card_is_needed);

    
endmodule