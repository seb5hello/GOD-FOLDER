`timescale 1ns / 1ps

/* 3-bit shift register */
module shift (
        // Clock (positive edge polarity)
        input clk,
        
        // Reset (active-high synchronous)
        input reset,
        
        // Input
        input in,
        
        // Output
        output [2:0] out
    );    
    
    // Add your logic here
    
endmodule