
module counter_ref(
    input clk,
    input reset,
    input tL,
    input tS,
    output trL,
    output trS,
    output hg,
    output hy,
    output hr,
    output fg,
    output fy,
    output fr);

    


endmodule