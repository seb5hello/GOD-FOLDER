module spi_parity_odd_fsm (
    input clk,
    input reset,
    input cs,
    input sample,
    input in,
    output parity_bit);

   
endmodule
