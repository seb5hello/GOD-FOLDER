module uart_retrans (
    input clk,
    input reset,
    input signal,
    input ack,
    output wire error,
    output wire [4:0] resend_count,
    output request_resend,
    output wire valid);

    
        
endmodule
