`timescale 1ns / 100ps

module seq_top (
    input  wire [0:0] clk,
    input  wire [0:0] reset,
    input  wire [0:0] update,
	input  wire [1:0] in,
	output reg  [0:0] p,
	output reg  [0:0] q
    );

endmodule
